`timescale 1ns / 1ps

module glitch_tube(

    );
endmodule
