`timescale 1ns / 1ps

//mode
//0: countdown
//1: winner each round
//2: final winner in scan_tube
//3: rejudge
module tube#(parameter mode=0)(
    input clk,
    input rst_n,
    output reg seg_out,
    output reg beep
);

   
    
    
endmodule